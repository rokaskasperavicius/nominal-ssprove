(** KEM-DEM example

  In this example, we follow the original SSP paper available at:
  https://eprint.iacr.org/2018/306

  In this file we first define the KEY pacakges and prove the single key lemma
  of the SSP paper. We then proceed to define the KEM-DEM packages and proving
  its security relative to that of the KEM and the DEM.
*)

Set Warnings "-notation-overridden,-ambiguous-paths,-notation-incompatible-format".
From mathcomp Require Import all_ssreflect all_algebra reals distr
  fingroup.fingroup realsum ssrnat ssreflect ssrfun ssrbool ssrnum eqtype choice
  seq.
Set Warnings "notation-overridden,ambiguous-paths,notation-incompatible-format".

From Crypt Require Import Axioms ChoiceAsOrd SubDistr Couplings
  UniformDistrLemmas FreeProbProg Theta_dens RulesStateProb UniformStateProb
  Package Prelude pkg_composition.

From Coq Require Import Utf8 Lia.
From extructures Require Import ord fset fmap.

From Equations Require Import Equations.
Require Equations.Prop.DepElim.

Set Equations With UIP.

Set Bullet Behavior "Strict Subproofs".
Set Default Goal Selector "!".
Set Primitive Projections.

Import Num.Def.
Import Num.Theory.
Import Order.POrderTheory.

Import PackageNotation.

From NominalSSP Require Import FsetSolve Nominal Fresh Pr NomPackage Disjoint.
Import FsetSolve.

#[local] Open Scope ring_scope.
#[local] Open Scope package_scope.

Section KEMDEM.

  (** We open a section in order to make local changes to global settings
      in the unlikely event that this module is imported somewhere else.
  *)
  Set Equations Transparent.

  (** In the SSP paper, bitstrings are used for the different data types.
      Instead we go for a more abstract types.
      In the cases where we need to be able to sample on these data types,
      we will first assume we have a (lossless) sub-distribution, and then
      define the types as the domain of these sub-distributions.
  *)

  (** Symmetric key *)
  Context (keyD : Op).
  Definition chKey := keyD.π1.

  (** Public and secret key *)
  Context (chPKey chSKey : choice_type).

  (** Plain text *)
  Context (chPlain : choice_type).

  (** We additionally require a "zero" in chPlain.

    Note that we don't require any structure on chPlain so this "zero" is only
    a "zero" in name a priori. Can be thought of as the 0 bitstring.
  *)
  Context (nullPlain : chPlain).

  (** Encrypted key

    This corresponds to the type of symmetric keys once encrypted.
  *)
  Context (ekeyD : Op).
  Definition chEKey := ekeyD.π1.

  (** Cipher text *)
  Context (cipherD : Op).
  Definition chCipher := cipherD.π1.

  (** Type notations *)

  Notation "'key" := (chKey) (in custom pack_type at level 2).
  Notation "'key" := (chKey) (at level 2) : package_scope.

  Notation "'pkey" := (chPKey) (in custom pack_type at level 2).
  Notation "'pkey" := (chPKey) (at level 2) : package_scope.

  Notation "'skey" := (chSKey) (in custom pack_type at level 2).
  Notation "'skey" := (chSKey) (at level 2) : package_scope.

  Notation "'plain" := (chPlain) (in custom pack_type at level 2).
  Notation "'plain" := (chPlain) (at level 2) : package_scope.

  Notation "'ekey" := (chEKey) (in custom pack_type at level 2).
  Notation "'ekey" := (chEKey) (at level 2) : package_scope.

  Notation "'cipher" := (chCipher) (in custom pack_type at level 2).
  Notation "'cipher" := (chCipher) (at level 2) : package_scope.

  (** Procedure names

    Under the hood, procedures are identified by natural numbers so we abstract
    them away by using distrinct coq-level identifiers.
  *)

  (* KEY *)
  Definition GEN := 0%N.
  Definition SET := 1%N.
  Definition GET := 2%N.

  (* KEM-CCA *)
  Definition KEMGEN := 6%N.
  Definition ENCAP := 7%N.
  Definition DECAP := 8%N.

  (* DEM-CCA *)
  Definition ENC := 9%N.
  Definition DEC := 10%N.

  (* PKE-CCA / MOD-CCA *)
  Definition PKGEN := 3%N.
  Definition PKENC := 4%N.
  Definition PKDEC := 5%N.

  (** Memory locations *)
  Definition k_loc : Location := ('option 'key ; 0%N).
  Definition pk_loc : Location := ('option 'pkey ; 1%N).
  Definition sk_loc : Location := ('option 'skey ; 2%N).
  Definition ek_loc : Location := ('option 'ekey ; 3%N).
  Definition c_loc : Location := ('option 'cipher ; 4%N).

  Definition pk_m_loc : Location := ('option 'pkey ; 5%N).
  Definition ek_m_loc : Location := ('option 'ekey ; 6%N).
  Definition c_m_loc : Location := ('option 'cipher ; 7%N).

  (** Some shorthands *)
  Definition IGEN := [interface #val #[ GEN ] : 'unit → 'unit ].
  Definition ISET := [interface #val #[ SET ] : 'key → 'unit ].
  Definition IGET := [interface #val #[GET] : 'unit → 'key ].

  (** PKE scheme

    A public-key encryption scheme comes with a key generation (a public and
    private key pair) and an encryption procedures (in the sense that they can
    use effects, typically sampling for the key generation procedure). It also
    comes with a pure (in particular deterministric) decryption function.
    The purity is denoted by the abscence of [code] in the return type.
  *)

  Record PKE_scheme := {
    PKE_kgen : code fset0 [interface] (chProd 'pkey 'skey) ;
    PKE_enc : 'pkey → 'plain → code fset0 [interface] (chProd 'ekey 'cipher) ;
    PKE_dec : 'skey → chProd 'ekey 'cipher → 'plain
  }.

  (** KEM scheme

    A key encapsulation mechanism comes with a key generation
    (public/private pair) and an encapsulation procedures as well as with a
    pure / deterministic decapsulation function.
  *)

  Record KEM_scheme := {
    KEM_kgen : code fset0 [interface] (chProd 'pkey 'skey) ;
    KEM_encap : 'pkey → code fset0 [interface] (chProd 'key 'ekey) ;
    KEM_decap : 'skey → 'ekey → 'key
  }.

  (** DEM scheme

    A data encapsulation mechanism comes with deterministric pure encryption
    and decryption functions. Both use a symmetric key.
  *)

  Record DEM_scheme := {
    DEM_enc : 'key → 'plain → 'cipher ;
    DEM_dec : 'key → 'cipher → 'plain
  }.

  (** We assume we are given a KEM and DEM schemes. *)
  Context (η : KEM_scheme).
  Context (θ : DEM_scheme).

  (** Specification of assumed schemes

    We assume the existence of a relation capturing which public key corresponds
    to which secret key. We furthermore require KEM_kgen to ensure that the
    keys it generates verify this relation.

    We use this relation to state the correctness of KEM_encap.

    The [⊢ₛ _ ⦃ _ ⦄] notation corresponds to unary specifications with only a
    post-condition on the result. They correspond to the diagonal of relational
    specifications, with the addition that state must be preserved.
  *)

  Context (pkey_pair : (chProd 'pkey 'skey) → Prop).
  Context (KEM_kgen_spec : ⊢ₛ η.(KEM_kgen) ⦃ pkey_pair ⦄).

  Definition encap_spec (pk : 'pkey) (kek : chProd 'key 'ekey) : Prop :=
    ∀ sk, pkey_pair (pk, sk) → η.(KEM_decap) sk kek.2 = kek.1.

  Context (KEM_encap_spec : ∀ pk, ⊢ₛ η.(KEM_encap) pk ⦃ encap_spec pk ⦄).

  (** KEY package *)

  (** The KEY package will only use one location: [k_loc] corresponding the
    stored key.
  *)
  Definition KEY_loc :=
    fset [:: k_loc ].

  (** Similarly, we define the export / output interface of the KEY package.

    The KEY package can generate a key [GEN] and then store its result in the
    location [k_loc] or alternatively it can set [SET] a key provided by the
    caller, finally in can return the stored key using [GET].
  *)
  Definition KEY_out :=
    [interface
      #val #[ GEN ] : 'unit → 'unit ;
      #val #[ SET ] : 'key → 'unit ;
      #val #[ GET ] : 'unit → 'key
    ].

  (** Definition of the KEY package *)
  Definition KEY : trimmed_package KEY_loc [interface] KEY_out :=
    [trimmed_package
      #def #[ GEN ] (_ : 'unit) : 'unit {
        k ← get k_loc ;;
        #assert (k == None) ;;
        k ← sample keyD ;;
        #put k_loc := Some k ;;
        @ret 'unit Datatypes.tt
      } ;
      #def #[ SET ] (k : 'key) : 'unit {
        k' ← get k_loc ;;
        #assert (k' == None) ;;
        #put k_loc := Some k ;;
        @ret 'unit Datatypes.tt
      } ;
      #def #[ GET ] (_ : 'unit) : 'key {
        k ← get k_loc ;;
        #assert (isSome k) as kSome ;;
        @ret 'key (getSome k kSome)
      }
    ].

  (** KEM package *)

  (** The KEM pacakge can refer to locations corresponding to a public and
    private asymetric keys, and to an encrypted symmetric key.
  *)
  Definition KEM_loc := fset [:: pk_loc ; sk_loc ; ek_loc ].

  (** The KEM packaee is parametrised by a boolean [b] depedning on which
    its import interface differs. If [b] is [true] it will be able to call
    the [SET] procedure, and if [b] is [false] it will be able to call the
    [GEN] one. In the paper [KEM true] corresponds to KEM⁰, while [KEM false]
    corresponds to KEM¹.
  *)
  Definition KEM_in b :=
    if b then ISET else IGEN.

  (** The KEM package will export a public and private key generation procedure
    [KEMGEM] that only returns the public one, an ecapsulation procedure [ENCAP]
    which will generate and encrypt a symmetric key, and a decpasulation
    procedure [DECAP] which returns a symmetric key given its encryption.
  *)
  Definition KEM_out :=
    [interface
      #val #[ KEMGEN ] : 'unit → 'pkey ;
      #val #[ ENCAP ] : 'unit → 'ekey ;
      #val #[ DECAP ] : 'ekey → 'key
    ].

  (** Here we add a hint to the [ssprove_valid_db] and [typeclass_instances]
    databases. The former database corresponds to what is used by the
    [ssprove_valid] tactic, while the latter corresponds to the built-in
    database used by type-class inference.
    This means that when Coq will have to prove the validity of a scheme, it
    will try to make use of the [valid_scheme] lemma that is a special case
    when the code does not import anything or use any state.
  *)
  Hint Extern 10 (ValidCode ?L ?I ?c.(prog)) =>
    eapply valid_scheme ; eapply c.(prog_valid)
    : typeclass_instances ssprove_valid_db.

  Definition KEM (b : bool) : trimmed_package KEM_loc (KEM_in b) KEM_out :=
    [trimmed_package
      #def #[ KEMGEN ] (_ : 'unit) : 'pkey {
        sk ← get sk_loc ;;
        #assert (sk == None) ;;
        '(pk, sk) ← η.(KEM_kgen) ;;
        #put pk_loc := Some pk ;;
        #put sk_loc := Some sk ;;
        @ret 'pkey pk
      } ;
      #def #[ ENCAP ] (_ : 'unit) : 'ekey {
        #import {sig #[ SET ] : 'key → 'unit } as SET ;;
        #import {sig #[ GEN ] : 'unit → 'unit } as GEN ;;
        pk ← get pk_loc ;;
        #assert (isSome pk) as pkSome ;;
        let pk := getSome pk pkSome in
        ek ← get ek_loc ;;
        #assert (ek == None) ;;
        '(k, ek) ← η.(KEM_encap) pk ;;
        #put ek_loc := Some ek ;;
        (if b then SET k else GEN Datatypes.tt) ;;
        ret ek
      } ;
      #def #[ DECAP ] (ek' : 'ekey) : 'key {
        sk ← get sk_loc ;;
        #assert (isSome sk) as skSome ;;
        let sk := getSome sk skSome in
        ek ← get ek_loc ;;
        #assert (ek != Some ek') ;;
        ret (η.(KEM_decap) sk ek')
      }
    ].

  (** KEM-CCA game

    The KEM-CCA game is obtained by composing the KEM and KEY packages, as well
    as the identity package. A game pair is described using a boolean-indexed
    function. Here, the only part that changes is the KEM package which is
    already indexed by a boolean.

    KEM-CCAᵇ = (KEMᵇ || ID) ∘ KEY
  *)

  Definition KEM_CCA_out :=
    [interface
      #val #[ KEMGEN ] : 'unit → 'pkey ;
      #val #[ ENCAP ] : 'unit → 'ekey ;
      #val #[ DECAP ] : 'ekey → 'key ;
      #val #[GET] : 'unit → 'key
    ].

  Definition KEM_CCA_loc :=
    KEM_loc :|: KEY_loc.

  (** Here we use Equations to generate a goal corresponding to the validity of
    the composed package as it is not inferred automatically.
    We call [ssprove_valid] which progresses as much as possible and then asks
    us to prove the remanining bits.

    Here and afterwards we use #[tactic=notac] to tell Equations not to
    preprocess the generated goals.
  *)
  Definition KEM_CCA b := dlink (dpar (KEM b) (nom_ID IGET)) KEY.

  #[local] Hint Unfold KEY_out IGET ISET IGEN : in_fset_eq.
  #[local] Hint Unfold KEM_in KEM_out KEM_CCA_out : in_fset_eq.

  Lemma idnts {n a b} : idents (fset (cons (n, a) b)) = n |: idents (fset b).
  Proof. 
    unfold idents.
    rewrite 2!imfset_fset //=.
    rewrite fset_cons //.
  Qed.
  Lemma idnts0 : idents fset0 = fset0.
  Proof. rewrite /idents imfset0 //. Qed.
  Lemma domm_emptym {T : ordType} {S : Type}
    : domm (@emptym T S) = fset0.
  Proof. unfold domm. simpl. rewrite fset0E //. Qed.
  #[local] Hint Rewrite domm_set @domm_ID @idnts @idnts0 @domm_emptym : in_fset_eq.

  #[export] Instance KEM_CCA_valid {b}
    : ValidPackage (loc (KEM_CCA b)) Game_import KEM_CCA_out (KEM_CCA b).
  Proof.
    unfold KEM_CCA.
    dprove_valid.
    destruct b; fset_solve.
  Qed.


  (** DEM package *)

  (** The DEM package only stores a cipher. *)
  Definition DEM_loc := fset [:: c_loc ].

  (** The DEM package can refer to the [GET] procedure. *)
  Definition DEM_in := IGET.

  (** The DEM package, produced from the DEM scheme θ, exports an encryption
    and a decryption procedures.
  *)
  Definition DEM_out :=
    [interface
      #val #[ ENC ] : 'plain → 'cipher ;
      #val #[ DEC ] : 'cipher → 'plain
    ].

  Definition DEM (b : bool) : trimmed_package DEM_loc DEM_in DEM_out :=
    [trimmed_package
      #def #[ ENC ] (m : 'plain) : 'cipher {
        #import {sig #[ GET ] : 'unit → 'key } as GET ;;
        c ← get c_loc ;;
        #assert (c == None) ;;
        k ← GET Datatypes.tt ;;
        let c := θ.(DEM_enc) k (if b then m else nullPlain) in
        #put c_loc := Some c ;;
        ret c
      } ;
      #def #[ DEC ] (c' : 'cipher) : 'plain {
        #import {sig #[ GET ] : 'unit → 'key } as GET ;;
        c ← get c_loc ;;
        #assert (c != Some c') ;;
        k ← GET Datatypes.tt ;;
        ret (θ.(DEM_dec) k c')
      }
    ].

  (** DEM-CCA game

    The DEM-CCA game is obtained by composing the DEM and KEY packages, as
    well as the indentity package.

    DEM-CCAᵇ = (DEMᵇ || ID) ∘ KEY
  *)

  Definition DEM_CCA_out :=
    [interface
      #val #[ GEN ] : 'unit → 'unit ;
      #val #[ ENC ] : 'plain → 'cipher ;
      #val #[ DEC ] : 'cipher → 'plain
    ].

  Definition DEM_CCA_loc :=
    DEM_loc :|: KEY_loc.

  Definition DEM_CCA b :=
    dlink (dpar (nom_ID IGEN) (DEM b)) KEY.

  #[local] Hint Unfold DEM_in DEM_out DEM_CCA_out : in_fset_eq.

  #[export] Instance DEM_CCA_valid {b}
    : ValidPackage (loc (DEM_CCA b)) Game_import DEM_CCA_out (DEM_CCA b).
  Proof.
    unfold DEM_CCA.
    dprove_valid.
  Qed.


  (** PKE-CCA *)

  Definition PKE_CCA_loc := fset [:: pk_loc ; sk_loc ; c_loc ; ek_loc ].

  Definition PKE_CCA_out :=
    [interface
      #val #[ PKGEN ] : 'unit → 'pkey ;
      #val #[ PKENC ] : 'plain → 'ekey × 'cipher ;
      #val #[ PKDEC ] : 'ekey × 'cipher → 'plain
    ].

  Definition PKE_CCA (ζ : PKE_scheme) b :
    trimmed_package PKE_CCA_loc Game_import PKE_CCA_out :=
    [trimmed_package
      #def #[ PKGEN ] (_ : 'unit) : 'pkey {
        sk ← get sk_loc ;;
        #assert (sk == None) ;;
        '(pk, sk) ← ζ.(PKE_kgen) ;;
        #put pk_loc := Some pk ;;
        #put sk_loc := Some sk ;;
        @ret 'pkey pk
      } ;
      #def #[ PKENC ] (m : 'plain) : 'ekey × 'cipher {
        pk ← get pk_loc ;;
        #assert (isSome pk) as pkSome ;;
        let pk := getSome pk pkSome in
        ek ← get ek_loc ;;
        #assert (ek == None) ;;
        c ← get c_loc ;;
        #assert (c == None) ;;
        '(ek, c) ← ζ.(PKE_enc) pk (if b then m else nullPlain) ;;
        #put ek_loc := Some ek ;;
        #put c_loc := Some c ;;
        @ret (chProd 'ekey 'cipher) (ek, c)
      } ;
      #def #[ PKDEC ] (c' : 'ekey × 'cipher) : 'plain {
        sk ← get sk_loc ;;
        #assert (isSome sk) as skSome ;;
        let sk := getSome sk skSome in
        ek ← get ek_loc ;;
        c ← get c_loc ;;
        #assert ((ek, c) != (Some c'.1, Some c'.2)) ;;
        ret (ζ.(PKE_dec) sk c')
      }
    ].

  (** MOD-CCA *)

  Definition MOD_CCA_loc :=
    fset [:: pk_m_loc ; c_m_loc ; ek_m_loc ].

  Definition MOD_CCA_in :=
    [interface
      #val #[ KEMGEN ] : 'unit → 'pkey ;
      #val #[ ENCAP ] : 'unit → 'ekey ;
      #val #[ DECAP ] : 'ekey → 'key ;
      #val #[ ENC ] : 'plain → 'cipher ;
      #val #[ DEC ] : 'cipher → 'plain
    ].

  Definition MOD_CCA_out :=
    PKE_CCA_out.

  Definition MOD_CCA (ζ : PKE_scheme) :
    trimmed_package MOD_CCA_loc MOD_CCA_in MOD_CCA_out :=
    [trimmed_package
      #def #[ PKGEN ] (_ : 'unit) : 'pkey {
        #import {sig #[ KEMGEN ] : 'unit → 'pkey } as KEMGEN ;;
        pk ← get pk_m_loc ;;
        #assert (pk == None) ;;
        pk ← KEMGEN Datatypes.tt ;;
        #put pk_m_loc := Some pk ;;
        ret pk
      } ;
      #def #[ PKENC ] (m : 'plain) : 'ekey × 'cipher {
        #import {sig #[ ENCAP ] : 'unit → 'ekey } as ENCAP ;;
        #import {sig #[ ENC ] : 'plain → 'cipher } as ENC ;;
        pk ← get pk_m_loc ;;
        #assert (isSome pk) ;;
        ek ← get ek_m_loc ;;
        #assert (ek == None) ;;
        c ← get c_m_loc ;;
        #assert (c ==  None) ;;
        ek ← ENCAP Datatypes.tt ;;
        #put ek_m_loc := Some ek ;;
        c ← ENC m ;;
        #put c_m_loc := Some c ;;
        @ret (chProd 'ekey 'cipher) (ek, c)
      } ;
      #def #[ PKDEC ] ('(ek', c') : 'ekey × 'cipher) : 'plain {
        #import {sig #[ DECAP ] : 'ekey → 'key } as DECAP ;;
        #import {sig #[ DEC ] : 'cipher → 'plain } as DEC ;;
        pk ← get pk_m_loc ;;
        #assert (isSome pk) ;;
        ek ← get ek_m_loc ;;
        c ← get c_m_loc ;;
        #assert ((ek, c) != (Some ek', Some c')) ;;
        if ek == Some ek'
        then (
          DEC c'
        )
        else (
          k' ← DECAP ek' ;;
          ret (θ.(DEM_dec) k' c')
        )
      }
    ].

  (** PKE scheme instance *)
  Definition KEM_DEM : PKE_scheme := {|
    PKE_kgen := η.(KEM_kgen) ;
    PKE_enc := λ pk m, {code
      '(k, ek) ← η.(KEM_encap) pk ;;
      let c := θ.(DEM_enc) k m in
      ret (ek, c)
    } ;
    PKE_dec := λ sk c,
      let '(ek, c) := c in
      let k := η.(KEM_decap) sk ek in
      θ.(DEM_dec) k c
  |}.

  (** Single key lemma *)

  (** Corresponds to Lemma 19.a in the SSP paper *)
  Lemma single_key_a :
    ∀ LD₀ LK₀ CK₀ CK₁ CD₀ CD₁ EK ED A,
      let K₀ := dlink (dpar CK₀ (nom_ID IGET)) KEY in
      let K₁ := dlink (dpar CK₁ (nom_ID IGET)) KEY in
      let D₀ := dlink (dpar (nom_ID IGEN) CD₀) KEY in
      let D₁ := dlink (dpar (nom_ID IGEN) CD₁) KEY in
      ValidPackage LD₀ IGET ED CD₀ →
      ValidPackage LD₀ IGET ED CD₁ →
      ValidPackage LK₀ ISET EK CK₀ →
      ValidPackage LK₀ IGEN EK CK₁ →
      Parable CK₀ (ID IGET) →
      Parable CK₁ (ID IGET) →
      Parable (ID IGEN) CD₀ →
      Parable (ID IGEN) CD₁ →
      trimmed ED CD₀ →
      trimmed ED CD₁ →
      trimmed EK CK₀ →
      trimmed EK CK₁ →
      AdvantageD (dlink (dpar CK₀ CD₀) KEY) (dlink (dpar CK₁ CD₁) KEY) A <=
      AdvantageD K₀ K₁ (dlink A (dpar (nom_ID EK) CD₀)) +
      AdvantageD D₀ D₁ (dlink A (dpar CK₁ (nom_ID ED))).
  Proof.
    intros LD₀ LK₀ CK₀ CK₁ CD₀ CD₁ EK ED A K₀ K₁ D₀ D₁.
    intros.
    advantage_trans (dlink (dpar CK₁ CD₀) KEY).
    erewrite -> (@AdvantageD_dpar_dlink_l _ _ _ _ _ _ _ _ _ (ISET :|: IGEN) IGET).
    (* why do we loop on first goal? with dprove_valid? *)
    2-10: try dprove_valid.
    erewrite -> (@AdvantageD_dpar_dlink_r _ _ _ _ _ _ _ _ _ IGEN IGET)
      ; dprove_valid.
  Qed.

  (** Corresponds to Lemma 19.b in the SSP paper *)
  Lemma single_key_b :
    ∀ LD₀ LK₀ CK₀ CK₁ CD₀ CD₁ EK ED A,
      let K₀ := dlink (dpar CK₀ (nom_ID IGET)) KEY in
      let K₁ := dlink (dpar CK₁ (nom_ID IGET)) KEY in
      let D₀ := dlink (dpar (nom_ID IGEN) CD₀) KEY in
      let D₁ := dlink (dpar (nom_ID IGEN) CD₁) KEY in
      ValidPackage LD₀ IGET ED CD₀ →
      ValidPackage LD₀ IGET ED CD₁ →
      ValidPackage LK₀ ISET EK CK₀ →
      ValidPackage LK₀ IGEN EK CK₁ →
      Parable CK₀ (ID IGET) →
      Parable CK₁ (ID IGET) →
      Parable (ID IGEN) CD₀ →
      Parable (ID IGEN) CD₁ →
      trimmed ED CD₀ →
      trimmed ED CD₁ →
      trimmed EK CK₀ →
      trimmed EK CK₁ →
      AdvantageD (dlink (dpar CK₀ CD₀) KEY) (dlink (dpar CK₀ CD₁) KEY) A <=
      AdvantageD K₀ K₁ (dlink A (dpar (nom_ID EK) CD₀)) +
      AdvantageD D₀ D₁ (dlink A (dpar CK₁ (nom_ID ED))) +
      AdvantageD K₀ K₁ (dlink A (dpar (nom_ID EK) CD₁)).
  Proof.
    intros LD₀ LK₀ CK₀ CK₁ CD₀ CD₁ EK ED A K₀ K₁ D₀ D₁.
    intros.
    advantage_trans (dlink (dpar CK₁ CD₁) KEY).
    eapply ler_add.
    - eapply single_key_a. all: eauto.
    (* De-idealising the core keying package *)
    - erewrite AdvantageD_sym.
      erewrite -> (@AdvantageD_dpar_dlink_l _ _ _ _ _ _ _ _ _ (ISET :|: IGEN) IGET)
        ; dprove_valid.
  Qed.

  (** Perfect indistinguishability with PKE-CCA

    We show that the package given by
    MOD_CCA KEM_DEM ∘ (KEM⁰ || DEMᵇ) ∘ KEY
    and which we call [Aux b], is perfectly indistinguishable from
    [PKE_CCA KEM_DEM b], which is the PKE-CCA game instantiated with the
    KEM-DEM instance we have.
  *)

  Definition Aux_loc :=
    MOD_CCA_loc :|: KEM_loc :|: DEM_loc :|: KEY_loc.

  Definition Aux b :=
    nom_link (MOD_CCA KEM_DEM) (nom_link (nom_par (KEM true) (DEM b)) KEY).

  #[local] Hint Unfold MOD_CCA_in : in_fset_eq.

  #[export] Instance Aux_valid {b : bool}
    : ValidPackage (loc (Aux b)) Game_import PKE_CCA_out (Aux b).
  Proof. unfold Aux. dprove_valid. Qed.

  Definition AuxD b :=
    dlink (MOD_CCA KEM_DEM) (dlink (dpar (KEM true) (DEM b)) KEY).

  #[export] Instance AuxD_valid {b}
    : ValidPackage (loc (AuxD b)) Game_import PKE_CCA_out (AuxD b).
  Proof.
    unfold AuxD.
    dprove_valid.
  Qed.

  (** We extend ssprove_code_simpl to use code_link_scheme.
    It says that linking a scheme with anything results in the scheme itself
    as a scheme does not import anything.
  *)
  Hint Extern 50 (_ = code_link _ _) =>
    rewrite code_link_scheme
    : ssprove_code_simpl.

  (** We extend swapping to schemes.
    This means that the ssprove_swap tactic will be able to swap any command
    with a scheme without asking a proof from the user.
  *)
  Hint Extern 40 (⊢ ⦃ _ ⦄ x ← ?s ;; y ← cmd _ ;; _ ≈ _ ⦃ _ ⦄) =>
    eapply r_swap_scheme_cmd ; ssprove_valid
    : ssprove_swap.

  (** Program equivalences

    In order to prove these equivalences, we will use an invariant that
    dismisses any changes made to the symmetric key location as it is only
    modified in one of the packages. This will be the [heap_ignore KEY_loc] bit
    in the following [inv] invariant.
    We need to extend this invariant with knowlegde about how the contents of
    some locations are related.
    With [triple_rhs pk_loc k_loc ek_loc PKE_inv] we say that the values
    corresponding to the public key, symmetric key and the encrypted symmetric
    key are always related by [PKE_inv] (described below).
    Similarly, [couple_lhs pk_loc sk_loc (sameSomeRel PkeyPair)] relates the
    public and secret keys by the relation [sameSomeRel PkeyPair]. It states
    that both must be [None], or both must be [Some pk] and [Some sk] such
    that [pk] and [sk] are related by [PkeyPair pk sk].
  *)

  (** This rephrasing of [pkey_pair] simply states that the stored public
    and private keys are indeed part of the same key pair, according to the
    specification of the KEM.
  *)
  Definition PkeyPair :=
    λ (pk : 'pkey) (sk : 'skey), pkey_pair (pk, sk).

  (** This states two things:
    - [k] and [ek] must both be set ([Some]) or unset ([None]);
    - whenever they are set, then the public key [pk] must as well and the three
    should be related by the functional specification [encap_spec] stating that
    [ek] is indeed the encryption of [k] using public key [pk].
  *)
  Definition PKE_inv (pk : 'option 'pkey) (k : 'option 'key) (ek : 'option 'ekey) :=
    match pk, k, ek with
    | Some pk, Some k, Some ek => encap_spec pk (k, ek)
    | Some pk, None, None => True
    | None, None, None => True
    | _, _, _ => False
    end.

  (*
  Definition derive_rhs (l l' : Location) (f : Value l.π1 → Value l'.π1) : precond :=
    couple_rhs l l' (λ a b, f a = b).

  Definition Derives_rhs (l l' : Location) f pre := Couples_rhs l l' (λ a b, f a = b) pre.
   *)

  Notation inv := (
    heap_ignore (MOD_CCA_loc :|: KEY_loc) ⋊
    couple_rhs pk_loc pk_m_loc eq ⋊
    couple_rhs ek_loc ek_m_loc eq ⋊
    couple_rhs c_loc c_m_loc eq ⋊
    triple_rhs pk_m_loc k_loc ek_loc PKE_inv ⋊
    couple_lhs pk_loc sk_loc (sameSomeRel PkeyPair)
  ).

  #[local]
  Hint Unfold PKE_CCA_loc MOD_CCA_loc Aux_loc : in_fset_eq.
  #[local]
  Hint Unfold KEM_loc DEM_loc KEY_loc : in_fset_eq.
  #[local]
  Hint Unfold Location : in_fset_eq.


  (** We have to show that [inv] is a valid invariant and while the
    [ssprove_invariant] does most of the work for us we still have some
    properties regarding the sets involved to prove
    (otherwise type inference would have solved it).
  *)
  Instance Invariant_inv {b} : Invariant PKE_CCA_loc (loc (Aux b)) inv.
  Proof.
    unfold Aux; simpl.
    ssprove_invariant; try done; fset_solve.
  Qed.

  (*
  Lemma Couples_rhs_Remembers_rhs {l l' v pre R} :
    Couples_rhs l l' R pre →
    (∀ v', R v v' → Remembers_rhs l' v' pre) →
    Remembers_rhs l v pre.
  Proof.
    intros cps rem s0 s1 preH.
    specialize (cps _ preH).
    unfold couple_rhs in cps.
    specialize (rem (get_heap s1 l')).
    unfold rem_rhs.
    specialize (rem _ _ _ _ preH).
   *)

  (*
     Search "r_rem".
  Search inv_conj.
  Lemma r_rem_suddenly_rhs :
    ∀ {A B : choiceType} (l : Location)
      (pre : precond) (c₀ : raw_code A) (c₁ : raw_code B) 
      (post : postcond A B),
        (∀ v, ⊢ ⦃ λ '(s₀, s₁), (pre ⋊ rem_rhs l v) (s₀, s₁) ⦄ c₀ ≈ c₁ ⦃ post ⦄)
          → ⊢ ⦃ λ '(s₀, s₁), pre (s₀, s₁) ⦄ c₀ ≈ c₁ ⦃ post ⦄.
  Proof.
    intros A B l pre c0 c1 post H.
    eapply rpre_weaken_rule. [ apply H |].
    intros s0 s1 preH.
    split; [ done |].
    reflexivity.
     Qed. *)


  (*
  Lemma r_rem_couple_rhs_cond:
    ∀ {A B : choiceType} (l l' : Location) (v : Value l.π1) 
      (R : Value l.π1 → Value l'.π1 → Prop) 
      (pre : precond) (c₀ : raw_code A) (c₁ : raw_code B) 
      (post : postcond A B),
      Couples_rhs l l' R pre
      → Remembers_rhs l v pre
          → (∀ v', ⊢ ⦃ λ '(s₀, s₁), (pre ⋊ rem_rhs l' v') (s₀, s₁) ⦄ c₀ ≈ c₁ ⦃ post ⦄)
            → ⊢ ⦃ λ '(s₀, s₁), pre (s₀, s₁) ⦄ c₀ ≈ c₁ ⦃ post ⦄.
  Proof.
    intros A B l l' v R pre c0 c1 post cps rem H.
    eapply rpre_weaken_rule.
    1: apply H.
    intros s0 s1 preH.
    (* 1: specialize (rem _ _ preH). *)
    simpl.
    split; [ done |].
    unfold rem_rhs.
    reflexivity.
    specialize (cps _ preH).
    specialize (rem _ _ preH).
    unfold couple_rhs in cps.
    unfold rem_rhs in rem.
    unfold rem_rhs.
    eapply r_rem_couple_rhs.
    

  Lemma Couples_rhs_Remembers_rhs {l l' v pre R} :
    Couples_rhs l l' R pre →
    Remembers_rhs l v pre →
    ∃ v', R v v' /\
    Remembers_rhs l' v' pre.
  Proof.
    intros cps rem.
    unfold Couples_rhs in cps.
    unfold Remembers_rhs in rem.
   *)

  Lemma r_get_vs_get_couples_rhs
     : ∀ {A B} (l l' : Location) (r₀ : Value l.π1 → raw_code A) 
         (r₁ : Value l'.π1 → raw_code B) (pre : precond) R
         (post : postcond A B),
         Syncs l pre →
         Couples_rhs l l' R pre →
         (∀ (x : Value l.π1) (x' : Value l'.π1), R x x' → ⊢ ⦃ λ '(s₀, s₁), (pre ⋊ rem_lhs l x ⋊ rem_rhs l' x') (s₀, s₁) ⦄
                 r₀ x ≈ r₁ x' ⦃ post ⦄) → ⊢ ⦃ λ '(s₀, s₁), pre (s₀, s₁) ⦄
              x ← get l ;;
              r₀ x ≈ x ← get l' ;;
                     r₁ x ⦃ post ⦄.
  Proof.
    intros A B l l' r₀ r₁ pre R post scs cps H.
    eapply r_get_remember_lhs => x.
    eapply r_get_remember_rhs => x'.
    eapply r_rem_couple_rhs.
    + do 2 apply Couples_rhs_conj_left; apply cps.
    + apply Remembers_rhs_from_tracked_lhs.
      2: by do 2 apply Syncs_conj.
      apply Remembers_lhs_conj_left, Remembers_lhs_conj_right.
      apply Remembers_lhs_rem_lhs.
    + apply Remembers_rhs_conj_right.
      apply Remembers_rhs_rem_rhs.
    + apply H.
  Qed.


  (** We show perfect equivalence in the general case where [b] stay abstract.
    This spares us the burden of proving roughly the same equivalence twice.
  *)
  Lemma PKE_CCA_perf :
    ∀ b, PKE_CCA KEM_DEM b ≈₀ Aux b.
  Proof.
    intro b.
    unfold Aux.
    (* We go to the relational logic with our invariant. *)
    eapply eq_rel_perf_ind with (inv := inv). 1: exact _.
    simplify_eq_rel m.
    (* rewrite !val_nom_link !val_nom_par /MOD_CCA /KEM /DEM /KEY !val_nom. *)
    all: ssprove_code_simpl.
    (* We are now in the realm of program logic *)
    - ssprove_code_simpl_more.
      ssprove_code_simpl.
      ssprove_swap_seq_rhs [:: 1 ; 0 ; 2 ; 1 ]%N.
      eapply r_get_vs_get_remember.
      1: ssprove_invariant; fset_solve. intro sk.
      ssprove_sync. intro skNone.
      eapply r_get_remember_rhs. intro pk.
      eapply (r_rem_couple_lhs pk_loc sk_loc). 1,3: exact _.
      1:{
        eapply Remembers_lhs_from_tracked_rhs.
        2: ssprove_invariant; fset_solve.
        intros s0 s1 [preH remH].
        do 6 move: preH => [preH _].
        move: preH => [_ preH].
        rewrite /rem_rhs preH remH //.
      }
      intro eps. destruct sk. 1: discriminate.
      destruct pk. 1: contradiction. simpl.
      eapply r_scheme_bind_spec. 1: eapply KEM_kgen_spec. intros [pk' sk'] pps.
      eapply r_put_vs_put.
      eapply r_put_vs_put.
      eapply r_put_rhs.
      ssprove_restore_mem.
      1:{
        ssprove_invariant; try auto.
        - intros s0 s1 hh.
          rewrite //= /heap_ignore.
          intros l H.
          rewrite (get_set_heap_neq _ pk_m_loc).
          2: fset_solve.
          destruct hh as [[[h _] h'] h''].
          simpl in h.
          destruct (l == sk_loc)%bool eqn:e.
          1: apply reflection_nonsense in e; subst; rewrite 2!get_set_heap_eq //.
          do 2 rewrite (get_set_heap_neq _ sk_loc) ?e //.
          destruct (l == pk_loc)%bool eqn:e'.
          1: apply reflection_nonsense in e'; subst; rewrite 2!get_set_heap_eq //.
          do 2 rewrite (get_set_heap_neq _ pk_loc) ?e' //.
          apply h, H.
        - intros s₀ s₁ hh. unfold triple_rhs in *. simpl in *.
          destruct hh as [[[hi ?] ?] e]. simpl in *.
          rewrite e in hi. get_heap_simpl.
          destruct (get_heap s₁ k_loc), (get_heap s₁ ek_loc).
          all: try contradiction.
          auto.
      }
      apply r_ret. auto.
    - ssprove_code_simpl_more.
      ssprove_code_simpl.
      ssprove_swap_seq_rhs [:: 5 ; 4 ; 3 ; 2 ; 1 ]%N.
      eapply r_get_remember_rhs => pk_m.
      eapply r_get_vs_get_remember. 1: ssprove_invariant; fset_solve. intro pk.
      eapply (r_rem_couple_rhs pk_loc pk_m_loc). 1,2,3: exact _.
      intros Eq; symmetry in Eq; subst.
      ssprove_sync. intro pkSome.
      destruct pk as [pk|]. 2: discriminate.
      simpl.
      ssprove_swap_seq_rhs [:: 3 ; 2 ; 1 ; 0 ]%N.
      eapply r_get_vs_get_remember. 1: ssprove_invariant; fset_solve. intro ek.
      eapply r_get_remind_rhs.
      1: {
        intros s0 s1 [[[[[[[[[_ H] _] _] _] _] _] _] _] H'].
        rewrite /rem_rhs -H H' //.
      }
      ssprove_sync. intro ekNone.
      rewrite ekNone. simpl.
      eapply r_get_vs_get_couples_rhs.
      1: ssprove_invariant; fset_solve.
      1: do 7 apply Couples_rhs_conj_left.
      1: apply Couples_rhs_conj_right.
      1: apply Couples_couple_rhs.
      intros c c' Eq; symmetry in Eq; subst.
      ssprove_sync. intro cNone.
      eapply r_scheme_bind_spec. 1: eapply KEM_encap_spec. intros [k' ek'] hkek.
      ssprove_code_simpl_more. ssprove_code_simpl.
      ssprove_code_simpl_more.
      ssprove_swap_seq_rhs [:: 3 ; 2 ; 1 ]%N.
      (* ssprove_contract_put_rhs. *)
      ssprove_swap_seq_rhs [:: 4 ; 3 ; 2 ; 1 ; 0 ]%N.
      eapply r_get_remind_rhs.
      1: apply Remembers_rhs_from_tracked_lhs.
      1: exact _.
      1: ssprove_invariant; fset_solve.
      rewrite cNone. simpl. ssprove_forget.
      ssprove_swap_seq_rhs [:: 1 ; 0 ]%N.
      eapply r_get_remember_rhs. intros k.
      eapply (r_rem_triple_rhs pk_m_loc k_loc ek_loc). 1-4: exact _. intro hpke.
      destruct ek. 1: discriminate.
      destruct k. 1: contradiction.
      simpl.
      ssprove_swap_seq_rhs [:: 1 ; 2 ; 0 ; 1 ]%N.
      ssprove_contract_put_get_rhs. simpl.
      apply r_put_rhs.
      apply r_put_vs_put.
      apply r_put_rhs.
      apply r_put_vs_put.
      apply r_put_rhs.
      ssprove_restore_mem.
      2: apply r_ret; auto.
      ssprove_invariant.
      2,3: reflexivity.
      1: rewrite -fset_cat.
      1: ssprove_invariant.
      intros s₀ s₁ hh. unfold triple_rhs in *. simpl in *.
      destruct hh as [[[[[[[hi epk] ?] ?] ?] ?] ?] ?]. simpl in *.
      get_heap_simpl.
      rewrite epk. simpl. auto.
    - destruct m as [ek' c']. simpl.
      ssprove_swap_seq_rhs [:: 1 ; 0 ; 2 ; 1 ]%N.
      ssprove_swap_seq_lhs [:: 1 ; 0 ; 2 ; 1 ]%N.
      eapply r_get_vs_get_couples_rhs.
      1: ssprove_invariant; fset_solve.
      1: exact _.
      intros ek ek_m Eq; symmetry in Eq; subst.
      eapply r_get_vs_get_couples_rhs.
      1: ssprove_invariant; fset_solve.
      1: exact _.
      intros c c_m Eq; symmetry in Eq; subst.
      eapply r_get_remember_rhs. intro pk.
      eapply r_get_remember_lhs. intro sk.
      eapply (r_rem_couple_lhs pk_loc sk_loc pk). 1,3: exact _.
      1: eapply Remembers_lhs_from_tracked_rhs.
      2: ssprove_invariant; fset_solve.
      1: {
        intros s0 s1 [[[[[[[[[[[_ H] _] _] _] _] _] _] _] _] H'] _].
        rewrite /rem_rhs H H' //.
      }

      intro eps.
      eapply sameSomeRel_sameSome in eps as eps'. rewrite eps'.
      ssprove_sync. intro skSome.
      ssprove_sync. intro neq.
      move: neq => /eqP neq.

      destruct (ek == Some ek')%bool eqn:eek.
      + move: eek => /eqP eek. subst ek.
        destruct (c != Some c') eqn:e.
        2:{ move: e => /eqP e. subst. contradiction. }
        rewrite eq_refl; simpl.
        eapply r_get_remind_rhs.
        1: eapply Remembers_rhs_from_tracked_lhs.
        1: exact _.
        1: ssprove_invariant; fset_solve.
        rewrite e.
        ssprove_code_simpl. simpl.
        ssprove_code_simpl. ssprove_code_simpl_more.
        eapply r_get_remember_rhs. intro k.
        eapply (r_rem_triple_rhs pk_m_loc k_loc ek_loc). 1,2,3: exact _.
        1: apply Remembers_rhs_from_tracked_lhs.
        1: exact _.
        1: ssprove_invariant; fset_solve.
        intro hpke.
        destruct sk as [sk|]. 2: discriminate.
        destruct pk as [pk|]. 2: contradiction.
        destruct k as [k|]. 2: contradiction.
        simpl. simpl in hpke. simpl in eps. unfold PkeyPair in eps.
        eapply hpke in eps as h. simpl in h. subst.
        ssprove_forget_all.
        apply r_ret. auto.
      + rewrite eek. ssprove_code_simpl_more.
        eapply r_get_remind_rhs.
        1: apply Remembers_rhs_from_tracked_lhs.
        1: exact _.
        1: ssprove_invariant; fset_solve.
        destruct sk as [sk|]. 2: discriminate.
        simpl.
        eapply r_get_remind_rhs.
        1: apply Remembers_rhs_from_tracked_lhs.
        1: exact _.
        1: ssprove_invariant; fset_solve.
        rewrite eek.
        simpl.
        ssprove_forget_all.
        apply r_ret; auto.
  Qed.


  (** Security theorem *)

  Lemma supp_trimmed_package {L I E} (P : trimmed_package L I E)
    : supp (trimmed_nom P) = supp L.
  Proof.
    done.
  Qed.

  Lemma supp1 {X : suppOrdType} {x : X} : supp (fset1 x) = supp x.
  Proof. apply fsetSupp1. Qed.

  (*
  #[local] Hint Rewrite @supp_fsetU : in_fset_eq.
  #[local] Hint Rewrite @fset_cons : in_fset_eq.
  #[local] Hint Rewrite @supp1 : in_fset_eq.
   *)

  Lemma supp_cons {X : suppOrdType} {x : X} {xs}
    : supp (fset (cons x xs)) = supp x :|: supp (fset xs).
  Proof. by rewrite fset_cons supp_fsetU supp1. Qed.

  Lemma supp_nil {X : suppOrdType}
    : supp (fset (@nil X)) = fset0.
  Proof. by rewrite -fset0E supp0. Qed.

  Lemma supp_Location (l : Location) : supp l = fset1 (atomize l.π2).
  Proof. destruct l. rewrite /supp //. Qed.

  #[local] Hint Rewrite @supp_cons @supp_nil @supp_Location : in_fset_eq.

  Lemma Aux_AuxD b : Aux b ≡ AuxD b.
  Proof.
    rewrite /Aux nom_link_dlink ?nom_link_dlink ?nom_par_dpar.
    1: reflexivity.
    1,2,3: rewrite /disj.
    2: rewrite s_nom_par.
    3: rewrite s_nom_link s_nom_par.
    1,2,3: rewrite !supp_trimmed_package.
    1,2,3: fset_solve.
  Qed.

  Theorem PKE_security :
    ∀ {LA} (A : nom_package),
      ValidPackage LA PKE_CCA_out A_export A →
      AdvantageP (PKE_CCA KEM_DEM) A <=
      AdvantageP KEM_CCA (dlink A
        (dlink (MOD_CCA KEM_DEM) (dpar (nom_ID KEM_out) (DEM true)))) +
      AdvantageP DEM_CCA (dlink A
        (dlink (MOD_CCA KEM_DEM) (dpar (KEM false) (nom_ID DEM_out)))) +
      AdvantageP KEM_CCA (dlink A
        (dlink (MOD_CCA KEM_DEM) (dpar (nom_ID KEM_out) (DEM false)))).
  Proof.
    intros LA A VA.
    unfold AdvantageP.
    erewrite (AdvantageD_perf_l (PKE_CCA_perf true)).
    erewrite (AdvantageD_perf_r (PKE_CCA_perf false)).
    rewrite 2!Aux_AuxD /AuxD.
    erewrite AdvantageD_dlink.
    eapply le_trans.
    + eapply (single_key_b _ _ _ (KEM false)).
      all: dprove_valid.
    + by erewrite dlink_assoc, dlink_assoc, dlink_assoc.
  Qed.
End KEMDEM.
